`define CLK_PERIOD 20.00ns

`ifndef BREAK_ERROR
  `define BREAK_ERROR 1
`endif

`ifndef TEST
  `define TEST 0
`endif


`ifndef TEST_FMA
  `define TEST_FMA 0
`endif

`ifndef TEST_SQRT
  `define TEST_SQRT 1
`endif
